module arithmetic_ops;
  int a=10, b=3;
  initial $display("a+b=%0d a*b=%0d a/b=%0d a%%b=%0d", a+b, a*b, a/b, a%b);
endmodule

