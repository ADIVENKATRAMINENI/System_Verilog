module if_else_basic;
  int x=10;
  initial if (x>5) $display("Greater than 5");
  else $display("Less or equal to 5");
endmodule

